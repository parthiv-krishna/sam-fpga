package instruction_decoder_params;
        localparam INPUT_SIGNAL_LENGTH = 32;
        localparam WRITE_DATA_LENGTH = 16;
        localparam WRITE_ADDRESS_LENGTH = 14;
	localparam READ_ADDRESS_LENGTH = 14;
endpackage
