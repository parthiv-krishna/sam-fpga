`timescale 1ns / 1ps

// instruction_decoder_tb: testbench for instruction_decoder

module instruction_decoder_tb(

    );
endmodule
